`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.04.2023 00:51:08
// Design Name: 
// Module Name: pc_4_adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//  This module isnt being used

/*module pc_4_adder(pc,pc4);

input [31:0] pc;
output reg [ 31:0] pc4;

always@(*)
begin
pc4 = pc + 4;
end

endmodule
*/
